* NGSPICE file created from OgueyAebischerBias.ext - technology: sky130A

.subckt nmos_5x a_408_100# a_n354_n158# a_n696_n100# a_n100_n158# a_n608_100# a_154_100#
+ a_408_n158# a_154_n158# a_n608_n158# a_n100_100# a_n354_100# VSUBS
X0 a_154_100# a_n696_n100# a_154_n158# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_n100_100# a_n696_n100# a_n100_n158# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_408_100# a_n696_n100# a_408_n158# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_n354_100# a_n696_n100# a_n354_n158# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_n608_100# a_n696_n100# a_n608_n158# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt pmos_7x a_408_100# a_662_100# a_n354_n158# a_n862_n158# w_n924_n194# a_n100_n158#
+ a_n960_n100# a_n608_100# a_n862_100# a_154_100# a_408_n158# a_154_n158# a_662_n158#
+ a_n608_n158# a_n100_100# a_n354_100#
X0 a_154_100# a_n960_n100# a_154_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_n100_100# a_n960_n100# a_n100_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_408_100# a_n960_n100# a_408_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_n862_100# a_n960_n100# a_n862_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_n354_100# a_n960_n100# a_n354_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X5 a_n608_100# a_n960_n100# a_n608_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 a_662_100# a_n960_n100# a_662_n158# w_n924_n194# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt OgueyAebischer_p7_n5 w_n44_400# pmos_7x_0/VSUBS m1_62_202# m1_220_n74# m1_n44_362#
+ m1_452_n204#
Xnmos_5x_1 m1_n44_362# m1_452_n204# m1_220_n74# pmos_7x_0/VSUBS m1_n44_362# m1_n44_362#
+ m1_452_n204# m1_452_n204# m1_452_n204# m1_220_n74# m1_n44_362# pmos_7x_0/VSUBS nmos_5x
Xpmos_7x_0 w_n44_400# w_n44_400# m1_220_n74# m1_62_202# w_n44_400# m1_n44_362# m1_n44_362#
+ w_n44_400# w_n44_400# w_n44_400# m1_220_n74# m1_220_n74# m1_62_202# m1_220_n74#
+ w_n44_400# w_n44_400# pmos_7x
.ends

.subckt nmos1x20_8x a_n354_2000# a_n862_2000# a_n100_2000# a_n950_n2000# a_408_n2058#
+ a_408_2000# a_916_2000# a_916_n2058# a_154_n2058# a_n100_n2058# a_662_n2058# a_154_2000#
+ a_n608_n2058# a_662_2000# a_n354_n2058# a_n608_2000# a_n862_n2058# VSUBS
X0 a_916_2000# a_n950_n2000# a_916_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X1 a_408_2000# a_n950_n2000# a_408_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X2 a_n608_2000# a_n950_n2000# a_n608_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X3 a_n100_2000# a_n950_n2000# a_n100_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X4 a_662_2000# a_n950_n2000# a_662_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X5 a_154_2000# a_n950_n2000# a_154_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X6 a_n862_2000# a_n950_n2000# a_n862_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X7 a_n354_2000# a_n950_n2000# a_n354_n2058# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt nmos_1x80_2x nmos1x20_8x_0/a_916_n2058# nmos1x20_8x_0/VSUBS nmos1x20_8x_0/a_662_n2058#
+ m1_n8_56# nmos1x20_8x_0/a_n608_n2058# nmos1x20_8x_0/a_n862_n2058#
Xnmos1x20_8x_0 m1_342_4064# m1_88_4064# m1_88_4064# m1_n8_56# m1_596_n154# m1_1358_4064#
+ m1_1104_4064# nmos1x20_8x_0/a_916_n2058# m1_850_n74# m1_850_n74# nmos1x20_8x_0/a_662_n2058#
+ m1_1104_4064# nmos1x20_8x_0/a_n608_n2058# m1_1358_4064# m1_596_n154# m1_342_4064#
+ nmos1x20_8x_0/a_n862_n2058# nmos1x20_8x_0/VSUBS nmos1x20_8x
.ends

.subckt OgueyAebischerBias vss vdd vbp vbn vbr vres
XOgueyAebischer_p7_n5_0 vdd vss vbr vbn vbp vres OgueyAebischer_p7_n5
Xnmos_1x80_2x_1 vss vss vss vbr vres vbr nmos_1x80_2x
.ends

