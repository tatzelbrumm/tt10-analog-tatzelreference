magic
tech sky130A
timestamp 1741712101
<< nwell >>
rect -362 240 145 364
<< poly >>
rect -233 287 -184 317
<< locali >>
rect -212 284 -195 320
<< metal1 >>
rect -215 181 -183 318
rect -167 221 -135 318
rect -44 -13 -14 281
rect 84 -13 114 281
<< via1 >>
rect -212 181 -186 207
rect -164 221 -138 247
rect -42 101 -16 127
rect 86 141 112 167
<< metal2 >>
rect -362 387 145 413
rect -362 221 145 247
rect -362 181 145 207
rect -362 141 145 167
rect -362 101 145 127
rect -362 61 145 87
rect -362 21 145 47
rect -362 -102 145 -76
rect -362 -142 145 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -281 0 1 302
box -81 -62 81 62
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 0 0 1 -34
box -163 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 0 0 1 302
box -163 -62 145 62
<< end >>
