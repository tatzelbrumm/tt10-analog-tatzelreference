magic
tech sky130A
magscale 1 2
timestamp 1741810117
<< nmos >>
rect -200 -831 200 769
<< ndiff >>
rect -258 757 -200 769
rect -258 -819 -246 757
rect -212 -819 -200 757
rect -258 -831 -200 -819
rect 200 757 258 769
rect 200 -819 212 757
rect 246 -819 258 757
rect 200 -831 258 -819
<< ndiffc >>
rect -246 -819 -212 757
rect 212 -819 246 757
<< poly >>
rect -200 841 200 857
rect -200 807 -184 841
rect 184 807 200 841
rect -200 769 200 807
rect -200 -857 200 -831
<< polycont >>
rect -184 807 184 841
<< locali >>
rect -200 807 -184 841
rect 184 807 200 841
rect -246 757 -212 773
rect -246 -835 -212 -819
rect 212 757 246 773
rect 212 -835 246 -819
<< viali >>
rect -184 807 184 841
rect -246 -819 -212 757
rect 212 -819 246 757
<< metal1 >>
rect -196 841 196 847
rect -196 807 -184 841
rect 184 807 196 841
rect -196 801 196 807
rect -252 757 -206 769
rect -252 -819 -246 757
rect -212 -819 -206 757
rect -252 -831 -206 -819
rect 206 757 252 769
rect 206 -819 212 757
rect 246 -819 252 757
rect 206 -831 252 -819
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
