magic
tech sky130A
timestamp 1741729423
use OgueyAebischer_p7_n5  OgueyAebischer_p7_n5_0
timestamp 1741324827
transform 1 0 0 0 1 0
box -22 -142 946 446
use ToBiasStartup  ToBiasStartup_0
timestamp 1741729423
transform 1 0 -166 0 1 0
box -367 -142 145 446
<< end >>
