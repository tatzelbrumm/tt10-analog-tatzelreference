magic
tech sky130A
timestamp 1741812120
<< nwell >>
rect -367 200 241 446
<< psubdiff >>
rect -20 -94 212 -92
rect -20 -111 -8 -94
rect 70 -111 122 -94
rect 200 -111 212 -94
rect -20 -113 212 -111
<< nsubdiff >>
rect -349 424 223 428
rect -349 407 -330 424
rect -242 407 -12 424
rect 204 407 223 424
rect -349 403 223 407
<< psubdiffcont >>
rect -8 -111 70 -94
rect 122 -111 200 -94
<< nsubdiffcont >>
rect -330 407 -242 424
rect -12 407 204 424
<< poly >>
rect -233 312 -184 317
rect -233 292 -212 312
rect -195 292 -184 312
rect -233 287 -184 292
<< polycont >>
rect -212 292 -195 312
<< locali >>
rect -338 407 -330 424
rect -242 407 -234 424
rect -20 407 -12 424
rect 204 407 212 424
rect -212 312 -195 320
rect -212 284 -195 292
rect -20 -111 -8 -94
rect 70 -111 122 -94
rect 200 -111 212 -94
<< viali >>
rect -330 407 -242 424
rect -12 407 76 424
rect 116 407 204 424
<< metal1 >>
rect -336 424 -236 428
rect -336 413 -330 424
rect -242 413 -236 424
rect -336 387 -333 413
rect -239 387 -236 413
rect -336 320 -236 387
rect -18 424 210 428
rect -18 413 -12 424
rect 76 413 116 424
rect 204 413 210 424
rect -18 387 -15 413
rect 79 403 113 413
rect 79 387 82 403
rect -18 320 82 387
rect 110 387 113 403
rect 207 387 210 413
rect 110 320 210 387
rect -268 247 -236 284
rect -268 221 -265 247
rect -239 221 -236 247
rect -215 207 -183 318
rect -71 247 -39 318
rect -71 221 -68 247
rect -42 221 -39 247
rect -215 181 -212 207
rect -186 181 -183 207
rect 52 127 82 281
rect 52 101 54 127
rect 80 101 82 127
rect -71 61 -68 87
rect -42 61 -39 87
rect -71 -37 -39 61
rect 52 0 82 101
rect 180 167 210 281
rect 180 141 182 167
rect 208 141 210 167
rect 180 0 210 141
rect -18 -116 82 -39
rect -18 -142 -15 -116
rect 79 -142 82 -116
rect 110 -116 210 -39
rect 110 -142 113 -116
rect 207 -142 210 -116
<< via1 >>
rect -333 407 -330 413
rect -330 407 -242 413
rect -242 407 -239 413
rect -333 387 -239 407
rect -15 407 -12 413
rect -12 407 76 413
rect 76 407 79 413
rect -15 387 79 407
rect 113 407 116 413
rect 116 407 204 413
rect 204 407 207 413
rect 113 387 207 407
rect -265 221 -239 247
rect -68 221 -42 247
rect -212 181 -186 207
rect 54 101 80 127
rect -68 61 -42 87
rect 182 141 208 167
rect -15 -142 79 -116
rect 113 -142 207 -116
<< metal2 >>
rect -367 387 -333 413
rect -239 387 -15 413
rect 79 387 113 413
rect 207 387 241 413
rect -268 221 -265 247
rect -239 221 -68 247
rect -42 221 -39 247
rect -367 181 -212 207
rect -186 181 241 207
rect -367 141 182 167
rect 208 141 241 167
rect -367 101 54 127
rect 80 101 241 127
rect -367 61 -68 87
rect -42 61 241 87
rect -367 -142 -15 -116
rect 79 -142 113 -116
rect 207 -142 241 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -286 0 1 302
box -81 -62 81 62
use nmos_8x2  nmos_8x2_0
timestamp 1741810117
transform -1 0 145 0 1 -2042
box 0 0 258 857
use nmos_8x2  nmos_8x2_1
timestamp 1741810117
transform -1 0 145 0 1 -1142
box 0 0 258 857
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 96 0 1 -21
box -163 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 96 0 1 302
box -163 -62 145 62
<< end >>
