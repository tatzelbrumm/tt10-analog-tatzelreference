magic
tech sky130A
timestamp 1741830316
<< nwell >>
rect -177 200 974 446
<< viali >>
rect 672 -203 760 -186
rect 799 -203 887 -186
<< metal1 >>
rect -144 101 -141 127
rect -115 101 -112 127
rect -144 -196 -112 101
rect -96 101 -93 127
rect 1 101 4 127
rect -96 -196 4 101
rect 909 101 912 127
rect 938 101 941 127
rect -144 -219 4 -196
rect -144 -2263 -112 -219
rect -96 -259 4 -219
rect 31 -102 34 -76
rect 128 -102 131 -76
rect 31 -259 131 -102
rect 666 -142 669 -116
rect 763 -142 766 -116
rect 666 -186 766 -142
rect 666 -203 672 -186
rect 760 -203 766 -186
rect 666 -259 766 -203
rect 793 -142 796 -116
rect 890 -142 893 -116
rect 793 -186 893 -142
rect 793 -203 799 -186
rect 887 -203 893 -186
rect 793 -259 893 -203
rect 909 -2263 941 101
<< via1 >>
rect -141 101 -115 127
rect -93 101 1 127
rect 912 101 938 127
rect 34 -102 128 -76
rect 669 -142 763 -116
rect 796 -142 890 -116
<< metal2 >>
rect -177 387 974 413
rect -177 181 974 207
rect -176 141 974 167
rect -177 101 -141 127
rect -115 101 -93 127
rect 1 101 912 127
rect 938 101 974 127
rect -177 -102 34 -76
rect 128 -102 974 -76
rect -177 -142 669 -116
rect 763 -142 796 -116
rect 890 -142 974 -116
use nmos_1x80_2x  nmos_1x80_2x_1
timestamp 1741828063
transform 1 0 -140 0 -1 -233
box -37 -77 1114 2135
use OgueyAebischer_p7_n5  OgueyAebischer_p7_n5_0
timestamp 1741829460
transform 1 0 0 0 1 0
box -22 -142 946 446
<< labels >>
rlabel metal2 -177 -142 -151 -116 1 vss
rlabel metal2 -177 387 -151 413 1 vdd
rlabel metal2 -177 181 -151 207 1 vbp
rlabel metal2 -176 141 -150 167 1 vbn
rlabel metal2 -177 101 -151 127 1 vbr
rlabel metal2 -177 -102 -151 -76 1 vres
<< end >>
