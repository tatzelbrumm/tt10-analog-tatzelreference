magic
tech sky130A
timestamp 1741834765
<< metal4 >>
rect 1503 22476 1533 22576
rect 1779 22476 1809 22576
rect 2055 22476 2085 22576
rect 2331 22476 2361 22576
rect 2607 22476 2637 22576
rect 2883 22476 2913 22576
rect 3159 22476 3189 22576
rect 3435 22476 3465 22576
rect 3711 22476 3741 22576
rect 3987 22476 4017 22576
rect 4263 22476 4293 22576
rect 4539 22476 4569 22576
rect 4815 22476 4845 22576
rect 5091 22476 5121 22576
rect 5367 22476 5397 22576
rect 5643 22476 5673 22576
rect 5919 22476 5949 22576
rect 6195 22476 6225 22576
rect 6471 22476 6501 22576
rect 6747 22476 6777 22576
rect 7023 22476 7053 22576
rect 7299 22476 7329 22576
rect 7575 22476 7605 22576
rect 7851 22476 7881 22576
rect 8127 22476 8157 22576
rect 8403 22476 8433 22576
rect 8679 22476 8709 22576
rect 8955 22476 8985 22576
rect 9231 22476 9261 22576
rect 9507 22476 9537 22576
rect 9783 22476 9813 22576
rect 10059 22476 10089 22576
rect 10335 22476 10365 22576
rect 10611 22476 10641 22576
rect 10887 22476 10917 22576
rect 11163 22476 11193 22576
rect 11439 22476 11469 22576
rect 11715 22476 11745 22576
rect 11991 22476 12021 22576
rect 12267 22476 12297 22576
rect 12543 22476 12573 22576
rect 12819 22476 12849 22576
rect 13095 22476 13125 22576
rect 100 500 300 22076
rect 400 500 600 22076
rect 700 500 900 22076
rect 93 0 183 100
rect 2025 0 2115 100
rect 3957 0 4047 100
rect 5889 0 5979 100
rect 7821 0 7911 100
rect 9753 0 9843 100
rect 11685 0 11775 100
rect 13617 0 13707 100
use tatzelreference_tile  tatzelreference_tile_0 ~/EDA/TinyTapeout/designs/tt10-analog-tatzelreference/mag
timestamp 1741834765
transform 1 0 0 0 1 0
box 0 0 14536 22576
<< labels >>
flabel metal4 s 12819 22476 12849 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 13095 22476 13125 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 12543 22476 12573 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 13617 0 13707 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 11685 0 11775 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 9753 0 9843 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 7821 0 7911 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 5889 0 5979 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 3957 0 4047 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 2025 0 2115 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 93 0 183 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 12267 22476 12297 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 11991 22476 12021 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 11715 22476 11745 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 11439 22476 11469 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 11163 22476 11193 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 10887 22476 10917 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 10611 22476 10641 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 10335 22476 10365 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 10059 22476 10089 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 9783 22476 9813 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 9507 22476 9537 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 9231 22476 9261 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 8955 22476 8985 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 8679 22476 8709 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 8403 22476 8433 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 8127 22476 8157 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 3435 22476 3465 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 3159 22476 3189 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 2883 22476 2913 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 2607 22476 2637 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 2331 22476 2361 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2055 22476 2085 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1779 22476 1809 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 1503 22476 1533 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 5643 22476 5673 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 5367 22476 5397 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 5091 22476 5121 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 4815 22476 4845 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 4539 22476 4569 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 4263 22476 4293 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 3987 22476 4017 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 3711 22476 3741 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 7851 22476 7881 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 7575 22476 7605 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 7299 22476 7329 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 7023 22476 7053 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 6747 22476 6777 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 6471 22476 6501 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 6195 22476 6225 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 5919 22476 5949 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 700 500 900 22076 1 FreeSans 200 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 14536 22576
<< end >>
