magic
tech sky130A
timestamp 1741330361
<< metal2 >>
rect -470 387 470 413
rect -470 181 470 207
rect -470 141 470 167
rect -470 101 470 127
rect -470 -102 470 -76
rect -470 -142 470 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -211 0 1 285
box -81 -62 81 62
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 0 0 1 3
box -127 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 0 0 1 285
box -145 -62 145 62
<< end >>
