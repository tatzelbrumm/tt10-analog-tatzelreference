magic
tech sky130A
timestamp 1740829677
<< nmos >>
rect 13 29 113 8029
<< ndiff >>
rect 13 8052 113 8058
rect 13 8035 19 8052
rect 107 8035 113 8052
rect 13 8029 113 8035
rect 13 23 113 29
rect 13 6 19 23
rect 107 6 113 23
rect 13 0 113 6
<< ndiffc >>
rect 19 8035 107 8052
rect 19 6 107 23
<< poly >>
rect 0 29 13 8029
rect 113 29 126 8029
<< locali >>
rect 11 8035 19 8052
rect 107 8035 115 8052
rect 11 6 19 23
rect 107 6 115 23
<< viali >>
rect 19 8035 107 8052
rect 19 6 107 23
<< metal1 >>
rect 13 8052 113 8055
rect 13 8035 19 8052
rect 107 8035 113 8052
rect 13 8032 113 8035
rect 13 23 113 26
rect 13 6 19 23
rect 107 6 113 23
rect 13 3 113 6
<< end >>
