magic
tech sky130A
timestamp 1741330361
<< metal2 >>
rect -292 387 145 413
rect -292 181 145 207
rect -292 141 145 167
rect -292 101 145 127
rect -292 -102 145 -76
rect -292 -142 145 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -211 0 1 285
box -81 -62 81 62
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 0 0 1 3
box -127 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 0 0 1 285
box -145 -62 145 62
<< end >>
