magic
tech sky130A
timestamp 1741351503
<< metal1 >>
rect -44 -13 -14 241
rect 84 -13 114 241
<< via1 >>
rect -42 101 -16 127
rect 86 141 112 167
<< metal2 >>
rect -292 387 145 413
rect -292 181 145 207
rect -292 141 145 167
rect -292 101 145 127
rect -292 61 145 87
rect -292 21 145 47
rect -292 -102 145 -76
rect -292 -142 145 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -211 0 1 262
box -81 -62 81 62
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 0 0 1 -34
box -127 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 0 0 1 262
box -145 -62 145 62
<< end >>
