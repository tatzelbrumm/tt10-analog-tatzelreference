magic
tech sky130A
timestamp 1741810884
<< nwell >>
rect -367 200 145 446
<< psubdiff >>
rect -116 -94 116 -92
rect -116 -111 -104 -94
rect -26 -111 26 -94
rect 104 -111 116 -94
rect -116 -113 116 -111
<< nsubdiff >>
rect -349 424 127 428
rect -349 407 -330 424
rect -242 407 -108 424
rect 108 407 127 424
rect -349 403 127 407
<< psubdiffcont >>
rect -104 -111 -26 -94
rect 26 -111 104 -94
<< nsubdiffcont >>
rect -330 407 -242 424
rect -108 407 108 424
<< poly >>
rect -233 312 -184 317
rect -233 292 -212 312
rect -195 292 -184 312
rect -233 287 -184 292
<< polycont >>
rect -212 292 -195 312
<< locali >>
rect -338 407 -330 424
rect -242 407 -234 424
rect -116 407 -108 424
rect 108 407 116 424
rect -212 312 -195 320
rect -212 284 -195 292
rect -116 -111 -104 -94
rect -26 -111 26 -94
rect 104 -111 116 -94
<< viali >>
rect -330 407 -242 424
rect -108 407 -20 424
rect 20 407 108 424
<< metal1 >>
rect -336 424 -236 428
rect -336 413 -330 424
rect -242 413 -236 424
rect -336 387 -333 413
rect -239 387 -236 413
rect -336 320 -236 387
rect -114 424 114 428
rect -114 413 -108 424
rect -20 413 20 424
rect 108 413 114 424
rect -114 387 -111 413
rect -17 403 17 413
rect -17 387 -14 403
rect -114 320 -14 387
rect 14 387 17 403
rect 111 387 114 413
rect 14 320 114 387
rect -268 247 -236 284
rect -268 221 -265 247
rect -239 221 -236 247
rect -215 207 -183 318
rect -167 247 -135 318
rect -167 221 -164 247
rect -138 221 -135 247
rect -215 181 -212 207
rect -186 181 -183 207
rect -44 127 -14 281
rect -44 101 -42 127
rect -16 101 -14 127
rect -167 61 -164 87
rect -138 61 -135 87
rect -167 -37 -135 61
rect -44 0 -14 101
rect 84 167 114 281
rect 84 141 86 167
rect 112 141 114 167
rect 84 0 114 141
rect -114 -116 -14 -39
rect -114 -142 -111 -116
rect -17 -142 -14 -116
rect 14 -116 114 -39
rect 14 -142 17 -116
rect 111 -142 114 -116
<< via1 >>
rect -333 407 -330 413
rect -330 407 -242 413
rect -242 407 -239 413
rect -333 387 -239 407
rect -111 407 -108 413
rect -108 407 -20 413
rect -20 407 -17 413
rect -111 387 -17 407
rect 17 407 20 413
rect 20 407 108 413
rect 108 407 111 413
rect 17 387 111 407
rect -265 221 -239 247
rect -164 221 -138 247
rect -212 181 -186 207
rect -42 101 -16 127
rect -164 61 -138 87
rect 86 141 112 167
rect -111 -142 -17 -116
rect 17 -142 111 -116
<< metal2 >>
rect -367 387 -333 413
rect -239 387 -111 413
rect -17 387 17 413
rect 111 387 145 413
rect -268 221 -265 247
rect -239 221 -164 247
rect -138 221 -135 247
rect -367 181 -212 207
rect -186 181 145 207
rect -367 141 86 167
rect 112 141 145 167
rect -367 101 -42 127
rect -16 101 145 127
rect -367 61 -164 87
rect -138 61 145 87
rect -367 -142 -111 -116
rect -17 -142 17 -116
rect 111 -142 145 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1740761609
transform 1 0 -286 0 1 302
box -81 -62 81 62
use nmos_8x2  nmos_8x2_0
timestamp 1741810117
transform -1 0 145 0 1 -2042
box 0 0 258 857
use nmos_8x2  nmos_8x2_1
timestamp 1741810117
transform -1 0 145 0 1 -1142
box 0 0 258 857
use shortnmos_2x  shortnmos_2x_0
timestamp 1740761609
transform 1 0 0 0 1 -21
box -163 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741318042
transform 1 0 0 0 1 302
box -163 -62 145 62
<< end >>
