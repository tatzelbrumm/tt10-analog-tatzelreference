magic
tech sky130A
timestamp 1741796374
<< psubdiff >>
rect -79 2085 1473 2106
rect -79 -49 1473 -28
<< locali >>
rect -79 2087 1473 2104
rect -79 -47 1473 -30
<< metal1 >>
rect 44 2109 47 2135
rect 141 2109 144 2135
rect 44 2032 144 2109
rect 425 2109 428 2135
rect 522 2109 525 2135
rect 171 2069 174 2095
rect 268 2069 271 2095
rect 171 2032 271 2069
rect 298 2069 301 2095
rect 395 2069 398 2095
rect 298 2032 398 2069
rect 425 2032 525 2109
rect 552 2109 555 2135
rect 649 2109 652 2135
rect 552 2032 652 2109
rect 933 2109 936 2135
rect 1030 2109 1033 2135
rect 679 2069 682 2095
rect 776 2069 779 2095
rect 679 2032 779 2069
rect 806 2069 809 2095
rect 903 2069 906 2095
rect 806 2032 906 2069
rect 933 2032 1033 2109
rect -4 28 28 2030
rect 1049 28 1081 2030
rect 298 -51 398 26
rect 425 -11 525 26
rect 425 -37 428 -11
rect 522 -37 525 -11
rect 552 -11 652 26
rect 552 -37 555 -11
rect 649 -37 652 -11
rect 298 -77 301 -51
rect 395 -77 398 -51
rect 679 -51 779 26
rect 679 -77 682 -51
rect 776 -77 779 -51
<< via1 >>
rect 47 2109 141 2135
rect 428 2109 522 2135
rect 174 2069 268 2095
rect 301 2069 395 2095
rect 555 2109 649 2135
rect 936 2109 1030 2135
rect 682 2069 776 2095
rect 809 2069 903 2095
rect 428 -37 522 -11
rect 555 -37 649 -11
rect 301 -77 395 -51
rect 682 -77 776 -51
<< metal2 >>
rect 44 2109 47 2135
rect 141 2109 428 2135
rect 522 2109 525 2135
rect 552 2109 555 2135
rect 649 2109 936 2135
rect 1030 2109 1033 2135
rect 171 2069 174 2095
rect 268 2069 301 2095
rect 395 2069 398 2095
rect 679 2069 682 2095
rect 776 2069 809 2095
rect 903 2069 906 2095
rect 425 -37 428 -11
rect 522 -37 555 -11
rect 649 -37 652 -11
rect 298 -77 301 -51
rect 395 -77 682 -51
rect 776 -77 779 -51
use nmos1x20_8x  nmos1x20_8x_0
timestamp 1741796374
transform 1 0 475 0 1 1029
box -475 -1029 603 1029
<< end >>
