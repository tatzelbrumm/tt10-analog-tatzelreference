magic
tech sky130A
timestamp 1741732016
<< error_s >>
rect 4437 1000 4537 1029
rect 4564 1000 4664 1029
rect 4691 1000 4791 1029
rect 4818 1000 4918 1029
rect 4945 1000 5045 1029
rect 5072 1000 5172 1029
rect 5199 1000 5299 1029
rect 5326 1000 5426 1029
<< isosubstrate >>
rect 0 0 14536 22576
<< metal4 >>
rect 11685 0 11775 200
rect 13617 0 13707 200
use OgueyAebischerBias  OgueyAebischerBias_0
timestamp 1741732016
transform 1 0 4533 0 1 3222
box -533 -2222 946 446
<< properties >>
string FIXED_BBOX 0 0 14536 22576
<< end >>
