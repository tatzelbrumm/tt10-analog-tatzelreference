magic
tech sky130A
timestamp 1741830316
use OgueyAebischerBias  OgueyAebischerBias_0
timestamp 1741830316
transform 1 0 0 0 1 0
box -177 -2368 974 446
use ToBiasStartup  ToBiasStartup_0
timestamp 1741828063
transform -1 0 -406 0 1 0
box -367 -2021 241 446
<< end >>
