magic
tech sky130A
<< nwell >>
rect -462 -97 462 97
<< pdiff >>
rect -431 -79 -331 79
rect -304 -79 -204 79
rect -177 -79 -77 79
rect -50 -79 50 79
rect 77 -79 177 79
rect 204 -79 304 79
rect 331 -79 431 79
<< pdiffc >>
rect -425 -73 -337 -56
rect -425 56 -337 73
rect -298 -73 -210 -56
rect -298 56 -210 73
rect -171 -73 -83 -56
rect -171 56 -83 73
rect -44 -73 44 -56
rect -44 56 44 73
rect 83 -73 171 -56
rect 83 56 171 73
rect 210 -73 298 -56
rect 210 56 298 73
rect 337 -73 425 -56
rect 337 56 425 73
<< poly >>
rect -454 -50 454 50
<< end >>
