magic
tech sky130A
magscale 1 2
timestamp 1741818438
<< error_s >>
rect -216 -4058 -158 -3205
rect 242 -4058 300 -3205
<< nwell >>
rect -734 400 482 892
<< psubdiff >>
rect -52 -188 412 -184
rect -52 -222 -28 -188
rect 128 -222 232 -188
rect 388 -222 412 -188
rect -52 -226 412 -222
<< nsubdiff >>
rect -698 848 434 856
rect -698 814 -660 848
rect -484 814 -36 848
rect 396 814 434 848
rect -698 806 434 814
<< psubdiffcont >>
rect -28 -222 128 -188
rect 232 -222 388 -188
<< nsubdiffcont >>
rect -660 814 -484 848
rect -36 814 396 848
<< poly >>
rect -466 624 -368 634
rect -466 584 -424 624
rect -390 584 -368 624
rect -466 574 -368 584
<< polycont >>
rect -424 584 -390 624
<< locali >>
rect -676 814 -660 848
rect -484 814 -468 848
rect -52 814 -36 848
rect 396 814 412 848
rect -424 624 -390 640
rect -424 568 -390 584
rect -52 -222 -28 -188
rect 128 -222 232 -188
rect 388 -222 412 -188
<< viali >>
rect -660 814 -484 848
rect -36 814 140 848
rect 220 814 396 848
<< metal1 >>
rect -672 848 -472 856
rect -672 826 -660 848
rect -484 826 -472 848
rect -48 848 408 856
rect -48 826 -36 848
rect 140 826 220 848
rect 396 826 408 848
rect -672 774 -666 826
rect -478 774 -472 826
rect -672 640 -472 774
rect -338 774 -332 826
rect -280 774 -274 826
rect -536 494 -472 568
rect -536 442 -530 494
rect -478 442 -472 494
rect -430 414 -366 636
rect -430 362 -424 414
rect -372 362 -366 414
rect -430 -532 -366 362
rect -338 -532 -274 774
rect -48 774 -42 826
rect 146 806 214 826
rect 146 774 152 806
rect -48 640 152 774
rect 208 774 214 806
rect 402 774 408 826
rect 208 640 408 774
rect -154 494 -90 636
rect -246 442 -240 494
rect -188 442 -182 494
rect -154 442 -148 494
rect -96 442 -90 494
rect -246 -532 -182 442
rect 92 254 152 562
rect 92 202 96 254
rect 148 202 152 254
rect -154 122 -148 174
rect -96 122 -90 174
rect -154 -532 -90 122
rect 92 0 152 202
rect 348 334 408 562
rect 348 282 352 334
rect 404 282 408 334
rect 348 0 408 282
rect -48 -232 152 -78
rect -48 -284 -42 -232
rect 146 -284 152 -232
rect 208 -232 408 -78
rect 208 -284 214 -232
rect 402 -284 408 -232
<< via1 >>
rect -666 814 -660 826
rect -660 814 -484 826
rect -484 814 -478 826
rect -666 774 -478 814
rect -332 774 -280 826
rect -530 442 -478 494
rect -424 362 -372 414
rect -42 814 -36 826
rect -36 814 140 826
rect 140 814 146 826
rect -42 774 146 814
rect 214 814 220 826
rect 220 814 396 826
rect 396 814 402 826
rect 214 774 402 814
rect -240 442 -188 494
rect -148 442 -96 494
rect 96 202 148 254
rect -148 122 -96 174
rect 352 282 404 334
rect -42 -284 146 -232
rect 214 -284 402 -232
<< metal2 >>
rect -734 774 -666 826
rect -478 774 -332 826
rect -280 774 -42 826
rect 146 774 214 826
rect 402 774 470 826
rect -536 442 -530 494
rect -478 442 -240 494
rect -188 442 -148 494
rect -96 442 -90 494
rect -734 362 -424 414
rect -372 362 470 414
rect -734 282 352 334
rect 404 282 470 334
rect -734 202 96 254
rect 148 202 470 254
rect -734 122 -148 174
rect -96 122 470 174
rect -734 -284 -42 -232
rect 146 -284 214 -232
rect 402 -284 470 -232
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1741818438
transform 1 0 -572 0 1 604
box -162 -124 162 124
use nmos_8x2  nmos_8x2_0
timestamp 1741818438
transform -1 0 300 0 1 -4084
box 0 0 516 1714
use nmos_8x2  nmos_8x2_1
timestamp 1741818438
transform -1 0 300 0 1 -2284
box 0 0 516 1714
use shortnmos_2x  shortnmos_2x_0
timestamp 1741818438
transform 1 0 180 0 1 -42
box -326 -88 254 88
use shortpmos_2x  shortpmos_2x_0
timestamp 1741818438
transform 1 0 180 0 1 604
box -326 -124 290 124
<< end >>
