magic
tech sky130A
timestamp 1741827447
use OgueyAebischerBias  OgueyAebischerBias_0
timestamp 1741827447
transform 1 0 0 0 1 0
box -177 -2368 974 446
use ToBiasStartup  ToBiasStartup_0
timestamp 1741827447
transform -1 0 -406 0 1 0
box -367 -2021 241 446
<< end >>
