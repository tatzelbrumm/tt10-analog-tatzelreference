magic
tech sky130A
timestamp 1741269935
<< error_s >>
rect 412 -114 512 -102
rect 415 -116 418 -114
rect 506 -116 509 -114
rect 412 -119 512 -116
rect 415 -128 509 -119
rect 412 -142 415 -139
rect 509 -142 512 -139
rect 415 -145 418 -142
rect 506 -145 509 -142
<< nwell >>
rect 0 392 924 446
<< psubdiff >>
rect 156 -94 768 -92
rect 156 -111 168 -94
rect 756 -111 768 -94
rect 156 -113 768 -111
<< nsubdiff >>
rect 18 424 906 428
rect 18 407 37 424
rect 886 407 906 424
rect 18 403 906 407
<< psubdiffcont >>
rect 168 -111 756 -94
<< nsubdiffcont >>
rect 37 407 886 424
<< locali >>
rect 29 407 37 424
rect 886 407 895 424
rect 29 353 895 370
rect 156 -111 168 -94
rect 756 -111 768 -94
<< viali >>
rect 418 -111 506 -94
<< metal1 >>
rect 31 373 131 428
rect 158 373 258 428
rect 285 373 385 428
rect 412 373 512 428
rect 539 373 639 428
rect 666 373 766 428
rect 793 373 893 428
rect 31 350 893 373
rect 99 127 131 244
rect 158 167 190 244
rect 158 141 161 167
rect 187 141 190 167
rect 226 181 229 207
rect 255 181 258 207
rect 99 101 102 127
rect 128 101 131 127
rect 226 67 258 181
rect 285 167 317 244
rect 412 207 444 244
rect 285 141 288 167
rect 314 141 317 167
rect 353 181 356 207
rect 382 181 385 207
rect 412 181 415 207
rect 441 181 444 207
rect 353 67 385 181
rect 539 167 571 244
rect 480 141 483 167
rect 509 141 512 167
rect 539 141 542 167
rect 568 141 571 167
rect 607 181 610 207
rect 636 181 639 207
rect 480 67 512 141
rect 607 67 639 181
rect 666 167 698 244
rect 666 141 669 167
rect 695 141 698 167
rect 734 181 737 207
rect 763 181 766 207
rect 734 67 766 181
rect 793 127 825 244
rect 793 101 796 127
rect 822 101 825 127
rect 226 -76 258 -39
rect 226 -102 229 -76
rect 255 -102 258 -76
rect 353 -76 385 -39
rect 353 -102 356 -76
rect 382 -102 385 -76
rect 412 -94 512 -39
rect 412 -111 418 -94
rect 506 -111 512 -94
rect 539 -76 571 -39
rect 539 -102 542 -76
rect 568 -102 571 -76
rect 666 -76 698 -39
rect 666 -102 669 -76
rect 695 -102 698 -76
rect 412 -114 512 -111
<< via1 >>
rect 161 141 187 167
rect 229 181 255 207
rect 102 101 128 127
rect 288 141 314 167
rect 356 181 382 207
rect 415 181 441 207
rect 483 141 509 167
rect 542 141 568 167
rect 610 181 636 207
rect 669 141 695 167
rect 737 181 763 207
rect 796 101 822 127
rect 229 -102 255 -76
rect 356 -102 382 -76
rect 542 -102 568 -76
rect 669 -102 695 -76
rect 415 -142 509 -116
<< metal2 >>
rect -9 181 229 207
rect 255 181 356 207
rect 382 181 415 207
rect 441 181 610 207
rect 636 181 737 207
rect 763 181 931 207
rect -9 141 161 167
rect 187 141 288 167
rect 314 141 483 167
rect 509 141 542 167
rect 568 141 669 167
rect 695 141 931 167
rect -9 101 102 127
rect 128 101 796 127
rect 822 101 931 127
rect -9 -102 229 -76
rect 255 -102 356 -76
rect 382 -102 542 -76
rect 568 -102 669 -76
rect 695 -102 931 -76
rect -9 -142 415 -116
rect 509 -142 931 -116
use nmos_5x  nmos_5x_1
timestamp 1740761609
transform -1 0 462 0 1 14
box -327 -79 327 79
use pmos_7x  pmos_7x_0
timestamp 1741269935
transform 1 0 462 0 1 297
box -462 -97 462 97
<< end >>
