magic
tech sky130A
timestamp 1741324827
<< nwell >>
rect 0 392 924 446
<< psubdiff >>
rect 156 -113 768 -92
<< nsubdiff >>
rect 18 403 906 428
<< psubdiffcont >>
rect 168 -111 756 -94
<< nsubdiffcont >>
rect 37 407 886 424
<< locali >>
rect 29 407 895 424
rect 29 353 895 370
rect 156 -111 768 -94
<< viali >>
rect 418 -111 506 -94
<< metal1 >>
rect 412 -142 512 -39
rect 226 -102 258 -39
rect 353 -102 385 -39
rect 539 -102 571 -39
rect 666 -102 698 -39
rect 31 350 893 373
rect 99 101 131 244
rect 158 141 190 244
rect 226 67 258 207
rect 285 141 317 244
rect 353 67 385 207
rect 412 181 444 244
rect 480 67 512 167
rect 539 141 571 244
rect 607 67 639 207
rect 666 141 698 244
rect 734 67 766 207
rect 793 101 825 244
rect 412 -114 512 -39
rect 31 350 131 428
rect 158 350 258 428
rect 285 350 385 428
rect 412 350 512 428
rect 539 350 639 428
rect 666 350 766 428
rect 793 350 893 428
<< via1 >>
rect 229 -102 255 -76
rect 356 -102 382 -76
rect 542 -102 568 -76
rect 669 -102 695 -76
rect 102 101 128 127
rect 161 141 187 167
rect 229 181 255 207
rect 288 141 314 167
rect 356 181 382 207
rect 415 181 441 207
rect 483 141 509 167
rect 542 141 568 167
rect 610 181 636 207
rect 669 141 695 167
rect 737 181 763 207
rect 796 101 822 127
rect 34 387 128 413
rect 161 387 255 413
rect 288 387 382 413
rect 415 387 509 413
rect 542 387 636 413
rect 669 387 763 413
rect 796 387 890 413
rect 415 -142 509 -116
<< metal2 >>
rect -9 -142 931 -116
rect -9 -102 931 -76
rect -9 181 931 207
rect -9 141 931 167
rect -9 101 931 127
rect -9 387 931 413
use nmos_5x  nmos_5x_1
timestamp 1740761609
transform -1 0 462 0 1 14
box -327 -79 327 79
use pmos_7x  pmos_7x_0
timestamp 1741324827
transform 1 0 462 0 1 297
box -462 -97 462 97
<< end >>
