magic
tech sky130A
timestamp 1740689597
<< comment >>
rect 0 0 14536 22576
<< properties >>
string FIXED_BBOX 0 0 14536 22576
<< end >>
