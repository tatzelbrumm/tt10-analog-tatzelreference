magic
tech sky130A
timestamp 1740761609
<< ndiff >>
rect -431 -1029 -331 1029
rect -304 -1029 -204 1029
rect -177 -1029 -77 1029
rect -50 -1029 50 1029
rect 77 -1029 177 1029
rect 204 -1029 304 1029
rect 331 -1029 431 1029
rect 331 -1029 431 1029
rect 458 -1029 558 1029
rect 458 -1029 558 1029
<< ndiffc >>
rect -425 -1023 -337 -1006
rect -425 1006 -337 1023
rect -298 -1023 -210 -1006
rect -298 1006 -210 1023
rect -171 -1023 -83 -1006
rect -171 1006 -83 1023
rect -44 -1023 44 -1006
rect -44 1006 44 1023
rect 83 -1023 171 -1006
rect 83 1006 171 1023
rect 210 -1023 298 -1006
rect 210 1006 298 1023
rect 337 -1023 425 -1006
rect 337 1006 425 1023
rect 464 -1023 552 -1006
rect 464 1006 552 1023
<< poly >>
rect -475 -1000 603 1000
<< polycont >>
rect -467 -995 -450 995
rect 577 -995 594 995
<< locali >>
rect -467 -1003 -450 1003
rect -433 -1023 -329 -1006
rect -433 1006 -329 1023
rect -306 -1023 -202 -1006
rect -306 1006 -202 1023
rect -179 -1023 -75 -1006
rect -179 1006 -75 1023
rect -52 -1023 52 -1006
rect -52 1006 52 1023
rect 75 -1023 179 -1006
rect 75 1006 179 1023
rect 202 -1023 306 -1006
rect 202 1006 306 1023
rect 329 -1023 433 -1006
rect 329 1006 433 1023
rect 456 -1023 560 -1006
rect 456 1006 560 1023
rect 577 -1003 594 1003
<< viali >>
rect -467 -995 -450 995
rect -425 -1023 -337 -1006
rect -425 1006 -337 1023
rect -298 -1023 -210 -1006
rect -298 1006 -210 1023
rect -171 -1023 -83 -1006
rect -171 1006 -83 1023
rect -44 -1023 44 -1006
rect -44 1006 44 1023
rect 83 -1023 171 -1006
rect 83 1006 171 1023
rect 210 -1023 298 -1006
rect 210 1006 298 1023
rect 337 -1023 425 -1006
rect 337 1006 425 1023
rect 464 -1023 552 -1006
rect 464 1006 552 1023
rect 577 -995 594 995
<< metal1 >>
rect -470 -1001 -447 1001
rect -431 -1026 -331 -1003
rect -431 1003 -331 1026
rect -304 -1026 -204 -1003
rect -304 1003 -204 1026
rect -177 -1026 -77 -1003
rect -177 1003 -77 1026
rect -50 -1026 50 -1003
rect -50 1003 50 1026
rect 77 -1026 177 -1003
rect 77 1003 177 1026
rect 204 -1026 304 -1003
rect 204 1003 304 1026
rect 331 -1026 431 -1003
rect 331 1003 431 1026
rect 458 -1026 558 -1003
rect 458 1003 558 1026
rect 574 -1001 597 1001
<< end >>
