magic
tech sky130A
timestamp 1741273084
use OgueyAebischer_p7_n5  OgueyAebischer_p7_n5_0
timestamp 1741273084
transform 1 0 0 0 1 0
box -9 -142 931 446
<< end >>
