magic
tech sky130A
timestamp 1740961960
<< metal2 >>
rect -9 181 931 207
rect -9 141 931 167
rect -9 101 931 127
<< end >>
