magic
tech sky130A
timestamp 1741827447
<< nwell >>
rect -367 200 241 446
<< psubdiff >>
rect -26 -94 206 -92
rect -26 -111 -14 -94
rect 64 -111 116 -94
rect 194 -111 206 -94
rect -26 -113 206 -111
rect -156 -186 198 -184
rect -156 -203 -137 -186
rect 179 -203 198 -186
rect -156 -205 198 -203
rect -156 -220 -135 -205
rect -156 -1077 -154 -220
rect -137 -1077 -135 -220
rect -156 -1092 -135 -1077
rect 177 -220 198 -205
rect 177 -1077 179 -220
rect 196 -1077 198 -220
rect 177 -1092 198 -1077
rect -156 -1094 198 -1092
rect -156 -1111 -137 -1094
rect 179 -1111 198 -1094
rect -156 -1113 198 -1111
rect -156 -1128 -135 -1113
rect -156 -1985 -154 -1128
rect -137 -1985 -135 -1128
rect -156 -2000 -135 -1985
rect 177 -1128 198 -1113
rect 177 -1985 179 -1128
rect 196 -1985 198 -1128
rect 177 -2000 198 -1985
rect -156 -2002 198 -2000
rect -156 -2019 -137 -2002
rect 179 -2019 198 -2002
rect -156 -2021 198 -2019
<< nsubdiff >>
rect -349 424 217 428
rect -349 407 -330 424
rect -242 407 -18 424
rect 198 407 217 424
rect -349 403 217 407
<< psubdiffcont >>
rect -14 -111 64 -94
rect 116 -111 194 -94
rect -137 -203 179 -186
rect -154 -1077 -137 -220
rect 179 -1077 196 -220
rect -137 -1111 179 -1094
rect -154 -1985 -137 -1128
rect 179 -1985 196 -1128
rect -137 -2019 179 -2002
<< nsubdiffcont >>
rect -330 407 -242 424
rect -18 407 198 424
<< poly >>
rect -236 312 -178 317
rect -236 292 -212 312
rect -186 292 -178 312
rect -236 287 -178 292
rect -82 312 -24 317
rect -82 292 -74 312
rect -48 292 -24 312
rect -82 287 -24 292
rect -128 -11 -24 -6
rect -128 -31 -120 -11
rect -94 -31 -24 -11
rect -128 -36 -24 -31
<< polycont >>
rect -212 292 -186 312
rect -74 292 -48 312
rect -120 -31 -94 -11
<< locali >>
rect -338 407 -330 424
rect -242 407 -234 424
rect -26 407 -18 424
rect 198 407 206 424
rect -212 312 -186 320
rect -212 284 -186 292
rect -74 312 -48 320
rect -74 284 -48 292
rect -120 -11 -94 -3
rect -120 -39 -94 -31
rect -26 -111 -14 -94
rect 64 -111 116 -94
rect 194 -111 206 -94
rect -154 -220 -137 -186
rect 179 -220 196 -186
rect -102 -1067 144 -263
rect -154 -1128 -137 -1077
rect 179 -1128 196 -1077
rect -103 -1975 143 -1171
rect -154 -2019 -137 -1985
rect 179 -2019 196 -1985
<< viali >>
rect -330 407 -242 424
rect -18 407 70 424
rect 110 407 198 424
rect -212 292 -186 312
rect -74 292 -48 312
rect -120 -31 -94 -11
<< metal1 >>
rect -336 424 -236 428
rect -336 413 -330 424
rect -242 413 -236 424
rect -24 424 204 428
rect -24 413 -18 424
rect 70 413 110 424
rect 198 413 204 424
rect -336 387 -333 413
rect -239 387 -236 413
rect -336 320 -236 387
rect -169 387 -166 413
rect -140 387 -137 413
rect -215 312 -183 318
rect -215 292 -212 312
rect -186 292 -183 312
rect -268 247 -236 284
rect -268 221 -265 247
rect -239 221 -236 247
rect -215 207 -183 292
rect -215 181 -212 207
rect -186 181 -183 207
rect -215 -1173 -183 181
rect -169 -1134 -137 387
rect -24 387 -21 413
rect 73 403 107 413
rect 73 387 76 403
rect -24 320 76 387
rect 104 387 107 403
rect 201 387 204 413
rect 104 320 204 387
rect -77 312 -45 318
rect -77 292 -74 312
rect -48 292 -45 312
rect -77 247 -45 292
rect -77 221 -74 247
rect -48 221 -45 247
rect -123 61 -120 87
rect -94 61 -91 87
rect -123 -11 -91 61
rect -123 -31 -120 -11
rect -94 -31 -91 -11
rect -123 -265 -91 -31
rect -77 -249 -45 221
rect 46 127 76 281
rect 46 101 48 127
rect 74 101 76 127
rect 46 0 76 101
rect 174 167 204 281
rect 174 141 176 167
rect 202 141 204 167
rect 174 0 204 141
rect -24 -116 76 -39
rect -24 -142 -21 -116
rect 73 -142 76 -116
rect 104 -116 204 -39
rect 104 -142 107 -116
rect 201 -142 204 -116
rect -123 -288 147 -265
rect -123 -1042 -91 -288
rect -123 -1065 147 -1042
rect -169 -1157 119 -1134
rect -215 -1196 147 -1173
rect -123 -1950 -91 -1196
rect -123 -1973 147 -1950
<< via1 >>
rect -333 407 -330 413
rect -330 407 -242 413
rect -242 407 -239 413
rect -333 387 -239 407
rect -166 387 -140 413
rect -265 221 -239 247
rect -212 181 -186 207
rect -21 407 -18 413
rect -18 407 70 413
rect 70 407 73 413
rect -21 387 73 407
rect 107 407 110 413
rect 110 407 198 413
rect 198 407 201 413
rect 107 387 201 407
rect -74 221 -48 247
rect -120 61 -94 87
rect 48 101 74 127
rect 176 141 202 167
rect -21 -142 73 -116
rect 107 -142 201 -116
<< metal2 >>
rect -367 387 -333 413
rect -239 387 -166 413
rect -140 387 -21 413
rect 73 387 107 413
rect 201 387 235 413
rect -268 221 -265 247
rect -239 221 -74 247
rect -48 221 -45 247
rect -367 181 -212 207
rect -186 181 235 207
rect -367 141 176 167
rect 202 141 235 167
rect -367 101 48 127
rect 74 101 235 127
rect -367 61 -120 87
rect -94 61 235 87
rect -367 -142 -21 -116
rect 73 -142 107 -116
rect 201 -142 235 -116
use flatpmos1x0.3  flatpmos1x0.3_0
timestamp 1741827447
transform 1 0 -286 0 1 302
box -81 -62 81 62
use nmos_8x2  nmos_8x2_0
timestamp 1741827447
transform -1 0 150 0 1 -1986
box 0 0 258 857
use nmos_8x2  nmos_8x2_1
timestamp 1741827447
transform -1 0 150 0 1 -1078
box 0 0 258 857
use shortnmos_2x  shortnmos_2x_0
timestamp 1741827447
transform 1 0 90 0 1 -21
box -127 -44 127 44
use shortpmos_2x  shortpmos_2x_0
timestamp 1741827447
transform 1 0 90 0 1 302
box -145 -62 145 62
<< end >>
