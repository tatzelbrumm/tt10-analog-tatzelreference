magic
tech sky130A
timestamp 1741833302
use OgueyAebischerBias  OgueyAebischerBias_0
timestamp 1741832991
transform 1 0 0 0 1 0
box -177 -2368 974 446
use ToBiasStartup  ToBiasStartup_0
timestamp 1741832991
transform -1 0 -406 0 1 0
box -367 -2021 235 446
<< labels >>
rlabel space -641 -142 -614 -116 1 vss
rlabel space -641 387 -614 413 1 vdd
rlabel space -641 181 -614 207 1 vbp
rlabel space -641 141 -614 167 1 vbn
rlabel space -641 101 -614 127 1 vbr
rlabel space -641 61 -614 87 1 disable
<< end >>
