magic
tech sky130A
timestamp 1740957648
<< locali >>
rect 29 353 895 370
<< metal1 >>
rect 31 350 893 373
rect 226 67 258 207
rect 353 67 385 207
rect 412 181 444 244
rect 607 67 639 207
rect 734 67 766 207
<< via1 >>
rect 229 181 255 207
rect 356 181 382 207
rect 415 181 441 207
rect 610 181 636 207
rect 737 181 763 207
<< metal2 >>
rect -9 181 931 207
rect -9 141 931 167
rect -9 101 931 127
use nmos_5x  nmos_5x_1
timestamp 1740957648
transform -1 0 462 0 1 14
box -327 -79 327 79
use pmos_7x  pmos_7x_0
timestamp 1740957648
transform 1 0 462 0 1 297
box -462 -97 462 97
<< end >>
