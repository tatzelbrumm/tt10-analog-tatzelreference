magic
tech sky130A
timestamp 1741829460
<< nwell >>
rect -22 200 946 446
<< psubdiff >>
rect 69 150 90 169
rect 69 -77 71 150
rect 88 -77 90 150
rect 69 -92 90 -77
rect 834 150 855 169
rect 834 -77 836 150
rect 853 -77 855 150
rect 834 -92 855 -77
rect 69 -94 855 -92
rect 69 -111 105 -94
rect 819 -111 855 -94
rect 69 -113 855 -111
<< nsubdiff >>
rect 18 424 906 428
rect 18 407 37 424
rect 886 407 906 424
rect 18 403 906 407
<< psubdiffcont >>
rect 71 -77 88 150
rect 836 -77 853 150
rect 105 -111 819 -94
<< nsubdiffcont >>
rect 37 407 886 424
<< locali >>
rect 29 407 37 424
rect 886 407 895 424
rect 29 353 895 370
rect 71 150 88 167
rect 71 -94 88 -77
rect 836 150 853 167
rect 836 -94 853 -77
rect 71 -111 105 -94
rect 819 -111 853 -94
<< viali >>
rect 418 -111 506 -94
<< metal1 >>
rect 31 413 131 428
rect 31 387 34 413
rect 128 387 131 413
rect 31 373 131 387
rect 158 413 258 428
rect 158 387 161 413
rect 255 387 258 413
rect 158 373 258 387
rect 285 413 385 428
rect 285 387 288 413
rect 382 387 385 413
rect 285 373 385 387
rect 412 413 512 428
rect 412 387 415 413
rect 509 387 512 413
rect 412 373 512 387
rect 539 413 639 428
rect 539 387 542 413
rect 636 387 639 413
rect 539 373 639 387
rect 666 413 766 428
rect 666 387 669 413
rect 763 387 766 413
rect 666 373 766 387
rect 793 413 893 428
rect 793 387 796 413
rect 890 387 893 413
rect 793 373 893 387
rect 31 350 893 373
rect -22 207 10 348
rect -22 181 -19 207
rect 7 181 10 207
rect 31 127 63 244
rect 158 167 190 244
rect 31 101 34 127
rect 60 101 63 127
rect 110 141 113 167
rect 139 141 142 167
rect 158 141 161 167
rect 187 141 190 167
rect 226 181 229 207
rect 255 181 258 207
rect 110 -37 142 141
rect 226 67 258 181
rect 285 167 317 244
rect 412 207 444 244
rect 285 141 288 167
rect 314 141 317 167
rect 353 181 356 207
rect 382 181 385 207
rect 412 181 415 207
rect 441 181 444 207
rect 353 67 385 181
rect 539 167 571 244
rect 480 141 483 167
rect 509 141 512 167
rect 539 141 542 167
rect 568 141 571 167
rect 607 181 610 207
rect 636 181 639 207
rect 480 67 512 141
rect 607 67 639 181
rect 666 167 698 244
rect 666 141 669 167
rect 695 141 698 167
rect 734 181 737 207
rect 763 181 766 207
rect 734 67 766 181
rect 782 141 785 167
rect 811 141 814 167
rect 782 -37 814 141
rect 861 127 893 244
rect 914 207 946 348
rect 914 181 917 207
rect 943 181 946 207
rect 861 101 864 127
rect 890 101 893 127
rect 226 -76 258 -39
rect 226 -102 229 -76
rect 255 -102 258 -76
rect 353 -76 385 -39
rect 353 -102 356 -76
rect 382 -102 385 -76
rect 412 -94 512 -39
rect 412 -111 418 -94
rect 506 -111 512 -94
rect 539 -76 571 -39
rect 539 -102 542 -76
rect 568 -102 571 -76
rect 666 -76 698 -39
rect 666 -102 669 -76
rect 695 -102 698 -76
rect 412 -116 512 -111
rect 412 -142 415 -116
rect 509 -142 512 -116
<< via1 >>
rect 34 387 128 413
rect 161 387 255 413
rect 288 387 382 413
rect 415 387 509 413
rect 542 387 636 413
rect 669 387 763 413
rect 796 387 890 413
rect -19 181 7 207
rect 34 101 60 127
rect 113 141 139 167
rect 161 141 187 167
rect 229 181 255 207
rect 288 141 314 167
rect 356 181 382 207
rect 415 181 441 207
rect 483 141 509 167
rect 542 141 568 167
rect 610 181 636 207
rect 669 141 695 167
rect 737 181 763 207
rect 785 141 811 167
rect 917 181 943 207
rect 864 101 890 127
rect 229 -102 255 -76
rect 356 -102 382 -76
rect 542 -102 568 -76
rect 669 -102 695 -76
rect 415 -142 509 -116
<< metal2 >>
rect -22 387 34 413
rect 128 387 161 413
rect 255 387 288 413
rect 382 387 415 413
rect 509 387 542 413
rect 636 387 669 413
rect 763 387 796 413
rect 890 387 946 413
rect -22 181 -19 207
rect 7 181 229 207
rect 255 181 356 207
rect 382 181 415 207
rect 441 181 610 207
rect 636 181 737 207
rect 763 181 917 207
rect 943 181 946 207
rect -22 141 113 167
rect 139 141 161 167
rect 187 141 288 167
rect 314 141 483 167
rect 509 141 542 167
rect 568 141 669 167
rect 695 141 785 167
rect 811 141 946 167
rect -22 101 34 127
rect 60 101 864 127
rect 890 101 946 127
rect -22 -102 229 -76
rect 255 -102 356 -76
rect 382 -102 542 -76
rect 568 -102 669 -76
rect 695 -102 946 -76
rect -22 -142 415 -116
rect 509 -142 946 -116
use nmos_5x  nmos_5x_1
timestamp 1741829076
transform -1 0 462 0 1 14
box -348 -79 348 79
use pmos_7x  pmos_7x_0
timestamp 1741829076
transform 1 0 462 0 1 297
box -480 -97 480 97
<< end >>
