magic
tech sky130A
timestamp 1740761609
<< ndiff >>
rect -431 -79 -331 79
rect -304 -79 -204 79
rect -177 -79 -77 79
rect -50 -79 50 79
rect 77 -79 177 79
rect 204 -79 304 79
rect 331 -79 431 79
<< ndiffc >>
rect -425 -73 -337 -56
rect -425 56 -337 73
rect -298 -73 -210 -56
rect -298 56 -210 73
rect -171 -73 -83 -56
rect -171 56 -83 73
rect -44 -73 44 -56
rect -44 56 44 73
rect 83 -73 171 -56
rect 83 56 171 73
rect 210 -73 298 -56
rect 210 56 298 73
rect 337 -73 425 -56
rect 337 56 425 73
<< poly >>
rect -454 -50 454 50
<< locali >>
rect -433 -73 -329 -56
rect -433 56 -329 73
rect -306 -73 -202 -56
rect -306 56 -202 73
rect -179 -73 -75 -56
rect -179 56 -75 73
rect -52 -73 52 -56
rect -52 56 52 73
rect 75 -73 179 -56
rect 75 56 179 73
rect 202 -73 306 -56
rect 202 56 306 73
rect 329 -73 433 -56
rect 329 56 433 73
<< viali >>
rect -425 -73 -337 -56
rect -425 56 -337 73
rect -298 -73 -210 -56
rect -298 56 -210 73
rect -171 -73 -83 -56
rect -171 56 -83 73
rect -44 -73 44 -56
rect -44 56 44 73
rect 83 -73 171 -56
rect 83 56 171 73
rect 210 -73 298 -56
rect 210 56 298 73
rect 337 -73 425 -56
rect 337 56 425 73
<< metal1 >>
rect -431 -76 -331 -53
rect -431 53 -331 76
rect -304 -76 -204 -53
rect -304 53 -204 76
rect -177 -76 -77 -53
rect -177 53 -77 76
rect -50 -76 50 -53
rect -50 53 50 76
rect 77 -76 177 -53
rect 77 53 177 76
rect 204 -76 304 -53
rect 204 53 304 76
rect 331 -76 431 -53
rect 331 53 431 76
<< end >>
