* NGSPICE file created from ToBiasStartup.ext - technology: sky130A

.subckt shortpmos_2x a_n254_n30# a_n228_n88# w_n290_n124# a_28_n88# a_n228_30#
X0 a_n228_30# a_n254_n30# a_n228_n88# w_n290_n124# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_n228_30# a_n254_n30# a_28_n88# w_n290_n124# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_BDGNGK a_200_n831# a_n200_n857# a_n258_n831# VSUBS
X0 a_200_n831# a_n200_n857# a_n258_n831# VSUBS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
.ends

.subckt nmos_8x2 sky130_fd_pr__nfet_01v8_BDGNGK_0/a_200_n831# sky130_fd_pr__nfet_01v8_BDGNGK_0/a_n200_n857#
+ sky130_fd_pr__nfet_01v8_BDGNGK_0/a_n258_n831# VSUBS
Xsky130_fd_pr__nfet_01v8_BDGNGK_0 sky130_fd_pr__nfet_01v8_BDGNGK_0/a_200_n831# sky130_fd_pr__nfet_01v8_BDGNGK_0/a_n200_n857#
+ sky130_fd_pr__nfet_01v8_BDGNGK_0/a_n258_n831# VSUBS sky130_fd_pr__nfet_01v8_BDGNGK
.ends

.subckt shortnmos_2x a_n254_n30# a_n228_n88# a_28_30# a_n228_30# VSUBS
X0 a_n228_30# a_n254_n30# a_n228_n88# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_28_30# a_n254_n30# a_n228_n88# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt flatpmos1x0.3 w_n162_n124# a_n100_n88# a_n126_n30# a_n100_30#
X0 a_n100_30# a_n126_n30# a_n100_n88# w_n162_n124# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt ToBiasStartup vss vdd vbp vbn vbr disable vkick
Xshortpmos_2x_0 vkick vbr vdd vbn vdd shortpmos_2x
Xnmos_8x2_0 vdd vbp vdd vss nmos_8x2
Xnmos_8x2_1 disable vkick disable vss nmos_8x2
Xshortnmos_2x_0 disable vss vbn vbr vss shortnmos_2x
Xflatpmos1x0.3_0 vdd vkick vbp vdd flatpmos1x0.3
.ends

