magic
tech sky130A
timestamp 1740829677
<< ndiff >>
rect 13 0 113 8058
<< ndiffc >>
rect 19 8035 107 8052
rect 19 6 107 23
<< poly >>
rect 0 29 126 8029
<< locali >>
rect 11 8035 115 8052
rect 11 6 115 23
<< viali >>
rect 19 8035 107 8052
rect 19 6 107 23
<< metal1 >>
rect 13 8032 113 8055
rect 13 3 113 26
<< end >>
